`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   02:13:48 01/04/2017
// Design Name:   top
// Module Name:   /home/mihailo/development/projects/layer_multiplex_nn/layer_multiplex_nn/tb_top.v
// Project Name:  layer_multiplex_nn
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: top
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb_forward;

    parameter LAYER_MAX       = 3,
              NUM_NEURON      = 7,              // max number of neurons
              INPUT_SIZE      = 9,              // width of the input signals
              WEIGHT_SIZE     = 17,             // width of the weight signals
              ADDR_SIZE       = 10,
              INPUT_FRACTION  = 8,              // number of bits below the radix point in the input
              WEIGHT_FRACTION = 8,              // number of bits below the radix point in the weight
              FRACTION_BITS   = 6;              // for the output of OUTPUT_SIZE, FRACTION_BITS is the number of bits 

    `include "../log2.v"

    reg [NUM_NEURON*NUM_NEURON*WEIGHT_SIZE-1:0] WEIGHTS [0:LAYER_MAX-1];

	// Inputs
	reg clk;
	reg rst;
	reg start;
	reg [NUM_NEURON*INPUT_SIZE-1:0] start_input;
    reg [NUM_NEURON*NUM_NEURON*WEIGHT_SIZE-1:0] weights;
    reg [log2(LAYER_MAX):0] layer_number;

	// Outputs
	wire [NUM_NEURON*INPUT_SIZE-1:0] final_output;
	wire final_output_valid;

    // Memories
    wire [9-1:0] output_mem [7-1:0];
    genvar i;
    generate
    for(i=0; i<7; i=i+1) begin: MEM
        assign output_mem[i] = final_output[i*9+:9];
    end
    endgenerate

	// Instantiate the Unit Under Test (UUT)
	forward #(
        .LAYER_MAX      (LAYER_MAX      ),
        .NUM_NEURON     (NUM_NEURON     ),
        .INPUT_SIZE     (INPUT_SIZE     ),
        .WEIGHT_SIZE    (WEIGHT_SIZE    ),
        .ADDR_SIZE      (ADDR_SIZE      ),
        .INPUT_FRACTION (INPUT_FRACTION ),
        .WEIGHT_FRACTION(WEIGHT_FRACTION),
        .FRACTION_BITS  (FRACTION_BITS  )
    ) uut (
		.clk(clk), 
		.rst(rst), 
		.start(start), 
        .weights(weights),
        .layer_number(layer_number),
		.start_input(start_input), 
		.final_output(final_output), 
		.final_output_valid(final_output_valid)
	);

    always
        #1 clk = ~clk;

	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 0;
		start = 0;
		start_input = 0;
        layer_number = 0;

        WEIGHTS[0] = 833'b11111111110010000000000000000000000000000101001100100000001100011001000000000000000000000000000000000011111111101110010111111111011100110000000001011100111111110101000110111111100111010110000000000000000000000000000000000000000000111111111111111110011100000000000101100101111111101111110001111110111101111100000000000000000000000000000000000000000001100101000000000010010010111111110010000110000000101100010000000001110100110000000000000000000000000000000000011111111100110110000000000000010100000000001001101111111110110010111111111100100001100000000000000000000000000000000000000000000100010101111111111111111111111111111100110000000001111101010000000100110101100000000000000000000000000000000001111111111010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000000;
        WEIGHTS[1] = 833'b00000000011000100111111110111000001111111100111110000000000110001100111111110010001000000000001110100100000000000111000111111111010001000000000101001000100000000110011100111111110001011110000000001111101011111111100010000000000000000111100000000010100000111111110111000010111111110011000010000000010100110011111111010110011000000001000011111111111111111110111111111110111110000000010001110010000000100010001111111111010111000000000000110010011111111111111100100000000000100011000000001000001101111111100110111011111111010101000000000000101010011111111101111010000000000011111001000000000000010111111111101110111100000000111011001000000010010011101111111101001010100000000110000110111111111010101010000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000000;
        WEIGHTS[2] = 833'b11111111001001100000000000111110111111111011110101011111111111010101111111110101011000000000000110111011111111111101000111111111101100111111111111001001111111111111001010111111111010101101111111110111101011111111100100011111111111110101000000000000011010111111111010111100000000000110101011111111101100101000000000001010010111111101111010101111111110111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000000;

        #20 rst = 1;
        #20 rst = 0;

        #20 start = 1;
            weights = WEIGHTS[0];
            layer_number = 0;
            start_input = 62'b010000010001011001000100011000000101000000000000000000011111111;
        #2  start = 0;

        #50 start = 1;
            weights = WEIGHTS[1];
            layer_number = 1;
        #2  start = 0;

        #50 start = 1;
            weights = WEIGHTS[2];
            layer_number = 1;
        #2  start = 0;


        // new input
        #100 start = 1;
            weights = WEIGHTS[0];
            layer_number = 0;
            start_input = 62'b010001100000111101001011110000011001000000000000000000011111111;
        #2  start = 0;

        #50 start = 1;
            weights = WEIGHTS[1];
            layer_number = 1;
        #2  start = 0;

        #50 start = 1;
            weights = WEIGHTS[2];
            layer_number = 1;
        #2  start = 0;


        // new input
        #100 start = 1;
            weights = WEIGHTS[0];
            layer_number = 0;
            start_input = 62'b010010111001001100010000010000101110000000000000000000011111111;
        #2  start = 0;

        #50 start = 1;
            weights = WEIGHTS[1];
            layer_number = 1;
        #2  start = 0;

        #50 start = 1;
            weights = WEIGHTS[2];
            layer_number = 1;
        #2  start = 0;

	end
      
endmodule

